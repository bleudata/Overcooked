//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Maya and Aarushi :)
// 
// Create Date: 11/14/2023
// Design Name: 
// Module Name: pickDropSprites.sv
// Project Name: Overcooked
// Target Devices: 
// Tool Versions: 
// Description: Bitmaps for the numbers 0 to 9 and : to display score and remaining time.
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module font_rom (input [8:0] addr, output [15:0] data);

    parameter ADDR_WIDTH = 9;
    parameter DATA_WIDTH = 16;
	logic [ADDR_WIDTH-1:0] addr_reg;
    parameter [0:351][DATA_WIDTH-1:0] ROM = {

// code x00
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00111111111100,
16'b00111111111100,
16'b11110000001111,
16'b11110000001111,
16'b11110000001111,
16'b11110000001111,
16'b11110000111111,
16'b11110000111111,
16'b11110011111111,
16'b11110011111111,
16'b11111111001111,
16'b11111111001111,
16'b11111100001111,
16'b11111100001111,
16'b11110000001111,
16'b11110000001111,
16'b11110000001111,
16'b11110000001111,
16'b00111111111100,
16'b00111111111100,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,

// code x01
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000011110000,
16'b00000011110000,
16'b00001111110000,
16'b00001111110000,
16'b00111111110000,
16'b00111111110000,
16'b00000011110000,
16'b00000011110000,
16'b00000011110000,
16'b00000011110000,
16'b00000011110000,
16'b00000011110000,
16'b00000011110000,
16'b00000011110000,
16'b00000011110000,
16'b00000011110000,
16'b00000011110000,
16'b00000011110000,
16'b00111111111111,
16'b00111111111111,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,

// code x02
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00111111111100,
16'b00111111111100,
16'b11110000001111,
16'b11110000001111,
16'b00000000001111,
16'b00000000001111,
16'b00000000111100,
16'b00000000111100,
16'b00000011110000,
16'b00000011110000,
16'b00001111000000,
16'b00001111000000,
16'b00111100000000,
16'b00111100000000,
16'b11110000000000,
16'b11110000000000,
16'b11110000001111,
16'b11110000001111,
16'b11111111111111,
16'b11111111111111,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,

// code x03
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00111111111100,
16'b00111111111100,
16'b11110000001111,
16'b11110000001111,
16'b00000000001111,
16'b00000000001111,
16'b00000000001111,
16'b00000000001111,
16'b00001111111100,
16'b00001111111100,
16'b00000000001111,
16'b00000000001111,
16'b00000000001111,
16'b00000000001111,
16'b00000000001111,
16'b00000000001111,
16'b11110000001111,
16'b11110000001111,
16'b00111111111100,
16'b00111111111100,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,

// code x04
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000111100,
16'b00000000111100,
16'b00000011111100,
16'b00000011111100,
16'b00001111111100,
16'b00001111111100,
16'b00111100111100,
16'b00111100111100,
16'b11110000111100,
16'b11110000111100,
16'b11111111111111,
16'b11111111111111,
16'b00000000111100,
16'b00000000111100,
16'b00000000111100,
16'b00000000111100,
16'b00000000111100,
16'b00000000111100,
16'b00000011111111,
16'b00000011111111,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,


// cod x05
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b11111111111111,
16'b11111111111111,
16'b11110000000000,
16'b11110000000000,
16'b11110000000000,
16'b11110000000000,
16'b11110000000000,
16'b11110000000000,
16'b11111111111100,
16'b11111111111100,
16'b00000000001111,
16'b00000000001111,
16'b00000000001111,
16'b00000000001111,
16'b00000000001111,
16'b00000000001111,
16'b11110000001111,
16'b11110000001111,
16'b00111111111100,
16'b00111111111100,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,


// code x06
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00001111110000,
16'b00001111110000,
16'b00111100000000,
16'b00111100000000,
16'b11110000000000,
16'b11110000000000,
16'b11110000000000,
16'b11110000000000,
16'b11111111111100,
16'b11111111111100,
16'b11110000001111,
16'b11110000001111,
16'b11110000001111,
16'b11110000001111,
16'b11110000001111,
16'b11110000001111,
16'b11110000001111,
16'b11110000001111,
16'b00111111111100,
16'b00111111111100,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,


// code x07
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b11111111111111,
16'b11111111111111,
16'b11110000001111,
16'b11110000001111,
16'b00000000001111,
16'b00000000001111,
16'b00000000001111,
16'b00000000001111,
16'b00000000111100,
16'b00000000111100,
16'b00000011110000,
16'b00000011110000,
16'b00001111000000,
16'b00001111000000,
16'b00001111000000,
16'b00001111000000,
16'b00001111000000,
16'b00001111000000,
16'b00001111000000,
16'b00001111000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,


// code x08
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00111111111100,
16'b00111111111100,
16'b11110000001111,
16'b11110000001111,
16'b11110000001111,
16'b11110000001111,
16'b11110000001111,
16'b11110000001111,
16'b00111111111100,
16'b00111111111100,
16'b11110000001111,
16'b11110000001111,
16'b11110000001111,
16'b11110000001111,
16'b11110000001111,
16'b11110000001111,
16'b11110000001111,
16'b11110000001111,
16'b00111111111100,
16'b00111111111100,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,

// code x09
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00111111111100,
16'b00111111111100,
16'b11110000001111,
16'b11110000001111,
16'b11110000001111,
16'b11110000001111,
16'b11110000001111,
16'b11110000001111,
16'b00111111111111,
16'b00111111111111,
16'b00000000001111,
16'b00000000001111,
16'b00000000001111,
16'b00000000001111,
16'b00000000001111,
16'b00000000001111,
16'b00000000111100,
16'b00000000111100,
16'b00111111110000,
16'b00111111110000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,

// code 0x0A
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000011110000,
16'b00000011110000,
16'b00000011110000,
16'b00000011110000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000011110000,
16'b00000011110000,
16'b00000011110000,
16'b00000011110000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000,
16'b00000000000000
};

	assign data = ROM[addr];

endmodule  